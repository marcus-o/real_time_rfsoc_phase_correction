`timescale 1ns / 1ps

module test();
  
    // instantiate bd
    test_bd_wrapper test_bd_i();

    initial begin

    end

endmodule